`define IMEM_FILE_TXT   "samples/fib_recursive.txt"
`define IMEM_FILE_MIF   "samples/fib_recursive.mif"

`define XBAR_MMIO_START 30'h0000
`define XBAR_MMIO_LIMIT 30'h03FF
`define XBAR_DATA_START 30'h0400
`define XBAR_DATA_LIMIT 30'h3FFF

`define XBAR_HEXD_ADDR0 30'h0008
