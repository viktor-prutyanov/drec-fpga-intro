/*
*   Replace with your clock divider
*/

module clk_div #(parameter X = 1)(
    input clk,

    output clk_out
);

endmodule
