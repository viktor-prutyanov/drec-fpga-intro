module alu(
    input [31:0]src_a,
    input [31:0]src_b,
    input [2:0]op,

    output reg [31:0]res
);

always @(*) begin
/*
* Problem 1:
* Write operations execution logic here.
*/
end

endmodule
