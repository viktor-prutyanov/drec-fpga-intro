/*
*   Replace with your hex display driver
*/

module hex_display(
    input clk,
    input [15:0]data,

    output [3:0]anodes,
    output [6:0]segments
);

endmodule
