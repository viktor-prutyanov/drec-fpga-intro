module top(
    input CLK
);

cpu_top cpu_top(.clk(CLK));

endmodule
