module counter #(parameter W = 16)(
    input clk,

    output [W - 1:0]q
);

/*
*   Write your code for counter of W bit width here
*/

endmodule
